`timescale 1ns/1ns

module tb_XOR_IO();

localparam WIDTH = 64;

logic 		[0:4][0:4][WIDTH-1:0] 	Xin;
logic 		[0:4][0:4][WIDTH-1:0] 	Xout;
logic 										X;

wire			[0:4][0:4][WIDTH-1:0] 	D;

XOR_IO XOR_IO_i(.*);

initial begin

	X = 0;

	Xin[0][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[1][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[2][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[3][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[4][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[0][1] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[1][1] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[2][1] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[3][1] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[4][1] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[0][2] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[1][2] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[2][2] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[3][2] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[4][2] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[0][3] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[1][3] = 64'hA3A3A3A3A3A3A3A3;	
	Xin[2][3] = 64'h0000000000000000;	
	Xin[3][3] = 64'h0000000000000000;	
	Xin[4][3] = 64'h0000000000000000;	
	Xin[0][4] = 64'h0000000000000000;	
	Xin[1][4] = 64'h0000000000000000;	
	Xin[2][4] = 64'h0000000000000000;	
	Xin[3][4] = 64'h0000000000000000;	
	Xin[4][4] = 64'h0000000000000000;
	
	Xout[0][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xout[1][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xout[2][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xout[3][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xout[4][0] = 64'hA3A3A3A3A3A3A3A3;	
	Xout[0][1] = 64'hA3A3A3A3A3A3A3A3;	
	Xout[1][1] = 64'hA3A3A3A3A3A3A3A3;	
	Xout[2][1] = 64'hA3A3A3A3A3A3A3A3;	
	Xout[3][1] = 64'h00000000000000C3;	
	Xout[4][1] = 64'h0000000000000000;	
	Xout[0][2] = 64'h0000000000000000;	
	Xout[1][2] = 64'h0000000000000000;	
	Xout[2][2] = 64'h0000000000000000;	
	Xout[3][2] = 64'h0000000000000000;	
	Xout[4][2] = 64'h0000000000000000;	
	Xout[0][3] = 64'h0000000000000000;	
	Xout[1][3] = 64'h8000000000000000;	
	Xout[2][3] = 64'h0000000000000000;	
	Xout[3][3] = 64'h0000000000000000;	
	Xout[4][3] = 64'h0000000000000000;	
	Xout[0][4] = 64'h0000000000000000;	
	Xout[1][4] = 64'h0000000000000000;	
	Xout[2][4] = 64'h0000000000000000;	
	Xout[3][4] = 64'h0000000000000000;	
	Xout[4][4] = 64'h0000000000000000;

	X = 1;
	
	#10 $stop;
	
end

endmodule 